* CPPSPICE - EXAMPLE 0 

L1 1 0 15e-2
I1 1 0 5
R1 1 2 10e3
C1 2 0 100e-6

*.OPTIONS SPARSE
.DC I1 0.0 10.0 1.0

.PLOT DC V(1) V(2)

*.TRAN 0.1 10

*.PLOT TRAN V(1) V(2)

*.AC LIN 100 0 1000

*.PLOT AC V(1) V(2)