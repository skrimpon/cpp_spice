L1 1 2 15e-2
V1 1 0 5 SIN (5 0.5 5 1 1 30)
R1 1 2 12e3
C1 2 0 100e-6

.tran 0.0001 3
.PLOT TRAN V(1) V(2)

.OPTIONS SPARSE METHOD = BE